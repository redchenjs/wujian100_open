/*
Copyright (c) 2019 Alibaba Group Holding Limited

Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

*/
module PAD_DIG_IO(
    OEN,
    IEN,
    OD,
    ID,
    PAD
);

input   OEN;
input   IEN;
output  ID;
input   OD;
inout   PAD;

// assign PAD = OEN ? 1'bz : OD;
// assign ID = IEN ? 1'bz : PAD;

IOBUF IOBUF_inst (
    .O(ID),         // Buffer output
    .IO(PAD),       // Buffer inout port (connect directly to top-level port)
    .I(OD),         // Buffer input
    .T(OEN &~ IEN)  // 3-state enable input, high=input, low=output
);

endmodule
